BZh91AY&SY!��m �߀Pxc����߰����`�=���d   m�I��X	D����I�4F@d4 z���쁥I&��       U??UT�h���&F �  JhA&�4�O"y  �a4�C���&L�20�&�db``
�"�S�b��Č�4 �=5��BH_*D�jH���^ζ톖���;^�.#�ImV�*%���]u��tj��I�DD		(  �   P �BQ�� �(
�iI��B��hK ��y�X@=G��N���`����ki�hR�*����gg�;qha$Z��LS�FB���N���f#&E��f.��A��oyO[��z�^�y���\����2-��V�B����׃V��+�n���4̐�z����|;�1����o��6[m�޸m��e����nm����s.&Sm���x�n[m�m��]̹m��m�m�ݶ�0�	w��ΐ���Cs��P����B�]e�&�<mpB){�DDD;�*�K��淋�������,K~O�uJ�Mݘ�n�-�;h[��R=��y�@:g�hM����{I($�b��1������*��/�Q1[>ļgQ������.w.k;v<.h��>p��>�	�� #E�^�W��/[)$�I/[ tЅ��|G�T@!�@6E $Fv��f{������pDQ l
U���<��UG��z������6��%FG���I$��<���JyH�]h$G=��@F&�����:���� a�D�Y4�`��|=��Rۉ�y:=Q��I$��4�R/����.x�-��R�]D��"�+%ΤR�E]����Żc�C]T�����j��DduxxGzI$�I%�����j�n�.{U�TNeV��Ɉ�z:�	�[<u\ݔ&#�"�Jq���w�G�G�7э$�I$���U~ed\�uTg��U2�x[��rGn�H�hGY���eQ;:vj����:X��w#�$�$��V���0���XX�呌����<�>�5�HF�kN|\Q'�I$���z��7�g���#
[�W��gN���3�%�$5��[�;G��9]��lړ�����I$�J���Nh�:��6`��C	����{��r�GDw��:mտ;z~���j�[y-�ń�»5�/d7��9
�Њ��!MHP���8;�*�K)e*�J�1ő�,�R�U*�R�e*�
U,���U*�S`�0�I�de��,M+5�T�K��L]՝�1f�=�ᶉg
X�k����ʳ�6{��@H;Nfj��<�F$��C�P�t�u�0ʐ��4�28z h
ilp&�Z��6����-��7�/��ʙ=%�b;���⽼�>!!��y{l�q%w���1(�>�obw���(�zR��n'V��O5�+5�7e�f�'��N����c��֘Տ%�m��f���=�eH��>Mϼ*S�O��P-��Hɰ�K@P��o�q��� �����nz)���$��V�p�j�AqƢb	"d$/
>���������p����_w�7��>r��=!��C��2Q�
�\&���I��ˁ�#j��.;S�N�1�L��1��j���h���� �h	�2Qr����<ņ��C�7W�E��������ߜ&%;��������;��(+�p�B
 ��̆����"�N�����f]�5yZ�:rmܚ�-�GD!�K8����#xB6m��h����+P��h����I��n&!����"�C;�WBʄ�������t�~.S]���p9��wm�M�Mb�r@t C��qw$S�	LF�